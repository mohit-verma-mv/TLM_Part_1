`include "uvm_macros.svh"
import uvm_pkg::*;

`include "seq_item.sv"

`include "driver.sv"
`include "converter.sv"
`include "stimulus.sv"

`include "producer.sv"
`include "consumer.sv"

`include "environment.sv"
`include "test.sv"

module top;
  
  initial
    begin
      run_test("test");
    end
  
endmodule